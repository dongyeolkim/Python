XPAD_AVDD1_0 TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDR_IN
XPAD_AVDD_3 TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDA_IN 
XPAD_AVDD_2 TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDA_IN 
XPAD_AVDD_1 TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDA_IN 
XPAD_AVDD_0 TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDA_IN 
XPAD_PLLVDD TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDPLL_IN 
XPAD_HVDD_2 TI1L1VDDIOK $PINS VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_HVDD_1 TI1L1VDDIOK $PINS VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_HVDD_0 TI1L1VDDIOK $PINS VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_SVDD_2 TI1L1XXAVDDNSUBK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN VDDNSUB=VDDS_IN 
XPAD_SVDD_1 TI1L1XXAVDDNSUBK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN VDDNSUB=VDDS_IN 
XPAD_SVDD_0 TI1L1XXAVDDNSUBK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN VDDNSUB=VDDS_IN 
XPAD_AVDD1_1 TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDR_IN
XPAD_DVDD_6 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_DVDD_5 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_DVDD_4 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_DVDD_3 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_DVDD_2 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_DVDD_1 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_DVDD_0 TI1L1VDDCOREK_DVDD_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_CVDD TI1L1AVDDEC33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVDD33OUT=VDDC_IN 
XPAD_HGND_2 TI1L1VSSK_HGND $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_HGND_1 TI1L1VSSK_HGND $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_HGND_0 TI1L1VSSK_HGND $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_AGND1 TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDR_IN 
XPAD_AGND_3 TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDA_IN
XPAD_AGND_2 TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDA_IN 
XPAD_AGND_1 TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDA_IN 
XPAD_AGND_0 TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDA_IN 
XPAD_DGND_5 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_DGND_4 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_DGND_3 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_DGND_2 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_DGND_1 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_DGND_0 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_CGND TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDC_IN 
XPAD_PLLGND TI1L1AVSS2DIECK2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN CVSSOUT=GNDPLL_IN 
XPAD_NCP TI1L1ABBOUT33K2_REV1 $PINS AVDD=VDDH_IN AVSS=GNDD_IN OUT=VREFN_PAD
XPAD_PCP TI1L1APPOUT33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN OUT=VREFP_PAD
XPAD_OSD TI1L1AIN33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN IN=OSD_PAD
XPAD_CN TI1L1AOUT33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN OUT=CN_PAD
XPAD_CP TI1L1AOUT33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN OUT=CP_PAD
XPAD_REXT TI1L1AOUT33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN OUT=REXT_PAD
XPAD_ISIN TI1L1AIN33K2 $PINS AVDD=VDDH_IN AVSS=GNDD_IN IN=ISIN_PAD
XPAD_DGND_6 TI1L1VSSK_DGND_PV2109K1 $PINS VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN 
XPAD_TE TI1L1IBN1CD1MEK $PINS IN=TE_PAD CFO=VDDH_IN OUT=w_te_pad_I IE=n_tie1_left 
+ VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN VSS3=GNDD_IN 
XPAD_CADDR TI1L1IBN1CD1MEK $PINS IN=CADDR_PAD CFO=VDDH_IN OUT=w_pad_chipaddr_I 
+ IE=n_tie1_left VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN VSS3=GNDD_IN 
XPAD_RSTB TI1L1IBN1CU1MEK $PINS IN=RSTB_PAD CFO=VDDH_IN OUT=w_rstb_pad_I 
+ IE=n_tie1_left VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN VSS3=GNDD_IN 
XPAD_STDBY TI1L1IBN1CD1MEK $PINS IN=STDBY_PAD CFO=VDDH_IN OUT=w_stdby_pad_I 
+ IE=n_tie1_left VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN VSS3=GNDD_IN 
XU_PAD_TIE_B tie_blk_v2 $PINS Z=por_out_I ZN=n_tie0_bot 
XU_PAD_TIE_T tie_blk_v2 $PINS Z=n_tie1_top ZN=n_tie0_top 
XU_PAD_TIE_R tie_blk_v2 $PINS Z=n_tie1_right ZN=n_tie0_right 
XU_PAD_TIE_L tie_blk_v2 $PINS Z=n_tie1_left ZN=n_tie0_left 
XPAD_X2 TI1L1XXP226OSC8N1K $PINS XCOM=xcom VDD=VDDD_IN VSS=GNDD_IN XO=X2_PAD 
+ CNT=osc_pad_ie_O CFO=VDDH_IN CHDRV=osc_drv_pad_O XOUT=mclk_pad_I VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_X1 TI1L1OSCXIK $PINS XI=X1_PAD XCOM=xcom VSS=GNDD_IN VDD=VDDD_IN VSS3=GNDD_IN VDD3=VDDH_IN
XU_buf_spidi_pad_I buf_blk_v1 $PINS A=w_spidi_pad_I Y=spidi_pad_I 
XU_buf_te_pad_I buf_blk_v1 $PINS A=w_te_pad_I Y=te_pad_I 
XU_buf_pad_chipaddr_I buf_blk_v1 $PINS A=w_pad_chipaddr_I Y=pad_chipaddr_I 
XU_buf_rstb_pad_I buf_blk_v1 $PINS A=w_rstb_pad_I Y=rstb_pad_I 
XU_buf_stdby_pad_I buf_blk_v1 $PINS A=w_stdby_pad_I Y=stdby_pad_I 
XPAD_MISO TI1L1IBN1CD1MEK $PINS IN=MISO_PAD CFO=VDDH_IN OUT=w_spidi_pad_I 
+ IE=spi_pad_ie_O VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN VSS3=GNDD_IN 
XPAD_LEDCTRL TI1L1ZBNC8S12ZSEK $PINS CHDRV=ledctrl_pad_drv_O IE=n_tie0_left 
+ VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN IO=LEDCTRL_PAD NOE=iv_ledctrl_pad_oen_O CFO=VDDH_IN 
+ IN=ledctrl_pad_O VSS3=GNDD_IN 
XPAD_PCLK TI1L1ZBNC8S12ZSEK $PINS CHDRV=pclk_drv_pad_O IE=n_tie0_right1 VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=PCLK_PAD NOE=iv_pclk_pad_oen_O CFO=VDDH_IN IN=isp_clk_pad_d_O VSS3=GNDD_IN 
XPAD_IRIS TI1L1ZBNC8S12ZSEK $PINS CHDRV=iris_pad_drv_O IE=n_tie0_right VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=IRIS_PAD NOE=iv_iris_pad_oen_O CFO=VDDH_IN IN=iris_pad_O VSS3=GNDD_IN 
XPAD_SDA TI1L1XXZNRBN1C6USU1MK_SDA $PINS NRST=VDDH_IN VDD=VDDD_IN VSS=GNDD_IN IO=SDA_PAD 
+ CFO=VDDH_IN OUT=sda_pad_I IN=iv_sda_pad_O IE=iv_sda_pad_O VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_SCL TI1L1XXZNRBN1C6USU1MK $PINS NRST=VDDH_IN VDD=VDDD_IN VSS=GNDD_IN IO=SCL_PAD 
+ CFO=VDDH_IN OUT=scl_pad_I IN=iv_scl_pad_O IE=n_tie1_right VSS3=GNDD_IN VDD3=VDDH_IN
XPAD_INT TI1L1ZBNC8S12ZSEK $PINS CHDRV=w1_int_pad_drv_O IE=n_tie0_top VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=INT_PAD NOE=iv_int_pad_oen_O CFO=VDDH_IN IN=w1_int_pad_O VSS3=GNDD_IN 
XU_w1_int_pad_drv_O buf_blk_v1 $PINS A=int_pad_drv_O Y=w1_int_pad_drv_O 
XU_w1_int_pad_O buf_blk_v1 $PINS A=int_pad_O Y=w1_int_pad_O 
XU_w1_vsync_pad_I buf_blk_v1 $PINS A=w1_vsync_pad_I Y=vsync_pad_I 
XU_w1_hsync_pad_ie_O buf_blk_v1 $PINS A=hsync_pad_ie_O Y=w1_hsync_pad_ie_O 
XU_w1_vsync_pad_ie_O buf_blk_v1 $PINS A=vsync_pad_ie_O Y=w1_vsync_pad_ie_O 
XPAD_CSB TI1L1ZBNC8S12ZSEK $PINS CHDRV=spi_pad_drv_O IE=n_tie0_left VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=CSB_PAD NOE=iv_spi_pad_oen_O CFO=VDDH_IN IN=spics_pad_O VSS3=GNDD_IN
XPAD_MOSI TI1L1ZBNC8S12ZSEK $PINS CHDRV=spi_pad_drv_O IE=n_tie0_left VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=MOSI_PAD NOE=iv_spido_pad_oen_O CFO=VDDH_IN IN=spido_pad_O VSS3=GNDD_IN
XPAD_SCK TI1L1ZBNC8S12ZSEK $PINS CHDRV=spi_pad_drv_O IE=n_tie0_left VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=SCK_PAD NOE=iv_spi_pad_oen_O CFO=VDDH_IN IN=spiclk_pad_O VSS3=GNDD_IN
XPAD_MIRS1 TI1L1ZBNC8S12ZSEK $PINS CHDRV=mirs_pad_drv_O IE=n_tie0_left VSS=GNDD_IN  
+ VDD=VDDD_IN VDD3=VDDH_IN IO=MIRS1_PAD NOE=iv_mirs_pad_oen_O CFO=VDDH_IN IN=mirs_pad_O[1] VSS3=GNDD_IN
XPAD_MIRS0 TI1L1ZBNC8S12ZSEK $PINS CHDRV=mirs_pad_drv_O IE=n_tie0_left VSS=GNDD_IN  
+ VDD=VDDD_IN VDD3=VDDH_IN IO=MIRS0_PAD NOE=iv_mirs_pad_oen_O CFO=VDDH_IN IN=mirs_pad_O[0] VSS3=GNDD_IN
XPAD_DC6 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_b_O IE=n_tie0_bot VSS=GNDD_IN  
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC6_PAD NOE=iv_dc6_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[6] VSS3=GNDD_IN
XPAD_DC7 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_b_O IE=dc7_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC7_PAD NOE=iv_dc7_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[10] 
+ IN=isp_data_smp_c_O[7] VSS3=GNDD_IN
XPAD_DC8 TI1L1ZBNC8S12USU1MEK $PINS CHDRV=pad_drv_b_O IE=dc8_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC8_PAD NOE=iv_dc8_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[0] 
+ IN=isp_data_smp_c_O[8] VSS3=GNDD_IN 
XPAD_DC9 TI1L1ZBNC8S12USU1MEK $PINS CHDRV=pad_drv_b_O IE=dc9_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC9_PAD NOE=iv_dc9_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[1] 
+ IN=isp_data_smp_c_O[9] VSS3=GNDD_IN 
XPAD_HSYNC TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=w1_pad_drv_t_O IE=w1_hsync_pad_ie_O 
+ VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN IO=HSYNC_PAD NOE=iv_hsync_pad_oen_O CFO=VDDH_IN 
+ OUT=w1_hsync_pad_I IN=hsync_smp_O VSS3=GNDD_IN 
XPAD_VSYNC TI1L1ZBNC8S12USU1MEK $PINS CHDRV=w1_pad_drv_t_O IE=w1_vsync_pad_ie_O 
+ VSS=GNDD_IN VDD=VDDD_IN VDD3=VDDH_IN IO=VSYNC_PAD NOE=iv_vsync_pad_oen_O CFO=VDDH_IN 
+ OUT=w1_vsync_pad_I IN=vsync_smp_O VSS3=GNDD_IN 
XU_w1_pad_drv_t_O buf_blk_v1 $PINS A=pad_drv_t_O Y=w1_pad_drv_t_O 
XU_w1_hsync_pad_I buf_blk_v1 $PINS A=w1_hsync_pad_I Y=hsync_pad_I 
XPAD_DY8 TI1L1ZBNC8S12USU1MEK $PINS CHDRV=pad_drv_r_O IE=dy8_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY8_PAD NOE=iv_dy8_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[8] 
+ IN=isp_data_smp_y_O[8] VSS3=GNDD_IN 
XPAD_DY9 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=dy9_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY9_PAD NOE=iv_dy9_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[9] 
+ IN=isp_data_smp_y_O[9] VSS3=GNDD_IN 
XPAD_DC0 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=n_tie0_right VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC0_PAD NOE=iv_dc0_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[0] VSS3=GNDD_IN 
XPAD_DC1 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=n_tie0_right VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC1_PAD NOE=iv_dc1_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[1] VSS3=GNDD_IN 
XPAD_DC2 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=n_tie0_right VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC2_PAD NOE=iv_dc2_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[2] VSS3=GNDD_IN 
XPAD_DC3 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=n_tie0_right VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC3_PAD NOE=iv_dc3_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[3] VSS3=GNDD_IN 
XPAD_DC4 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=n_tie0_right VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC4_PAD NOE=iv_dc4_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[4] VSS3=GNDD_IN 
XPAD_DC5 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_b_O IE=n_tie0_bot VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DC5_PAD NOE=iv_dc5_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_c_O[5] VSS3=GNDD_IN 
XPAD_DY0 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_t_O IE=n_tie0_top VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY0_PAD NOE=iv_motion_pad_oen_O CFO=VDDH_IN 
+ IN=isp_data_smp_y_O[0] VSS3=GNDD_IN 
XPAD_DY1 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_t_O IE=n_tie0_top VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY1_PAD NOE=iv_dy1_pad_oen_O CFO=VDDH_IN IN=isp_data_smp_y_O[1] VSS3=GNDD_IN 
XPAD_DY2 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_t_O IE=dy2_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY2_PAD NOE=iv_dy2_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[2] 
+ IN=isp_data_smp_y_O[2] VSS3=GNDD_IN 
XPAD_DY3 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_t_O IE=dy3_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY3_PAD NOE=iv_dy3_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[3] 
+ IN=isp_data_smp_y_O[3] VSS3=GNDD_IN 
XPAD_DY4 TI1L1ZBNC8S12USU1MEK $PINS CHDRV=pad_drv_t_O IE=dy4_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY4_PAD NOE=iv_dy4_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[4] 
+ IN=isp_data_smp_y_O[4] VSS3=GNDD_IN 
XPAD_DY5 TI1L1ZBNC8S12USU1MEK $PINS CHDRV=pad_drv_t_O IE=dy5_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY5_PAD NOE=iv_dy5_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[5] 
+ IN=isp_data_smp_y_O[5] VSS3=GNDD_IN 
XPAD_DY6 TI1L1ZBNC8S12USU1MEK $PINS CHDRV=pad_drv_r_O IE=dy6_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY6_PAD NOE=iv_dy6_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[6] 
+ IN=isp_data_smp_y_O[6] VSS3=GNDD_IN 
XPAD_DY7 TI1L1ZBNC8S12DSD1MEK $PINS CHDRV=pad_drv_r_O IE=dy7_pad_ie_O VSS=GNDD_IN 
+ VDD=VDDD_IN VDD3=VDDH_IN IO=DY7_PAD NOE=iv_dy7_pad_oen_O CFO=VDDH_IN OUT=scan_in_pad_I[7] 
+ IN=isp_data_smp_y_O[7] VSS3=GNDD_IN  
XU_PAD_TIE_R1 tie_blk_v2 $PINS ZN=n_tie0_right1 
Xana_filler_133 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_153 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_306 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_307 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_308 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_309 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_1 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_2 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_3 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_4 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_5 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_6 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_7 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_8 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_9 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_10 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_11 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_12 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_22 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_24 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_25 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_26 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_27 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_30 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_31 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_35 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_37 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_38 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_41 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_42 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_43 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_44 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_45 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_46 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_47 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_49 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_50 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_52 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_53 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_54 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_55 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_301 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_58 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_59 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_61 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_62 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_63 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_64 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_304 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_67 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_68 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_70 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_71 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_72 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_73 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_75 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_76 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_77 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_79 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_80 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_82 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_83 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_84 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_85 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_86 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_87 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_305 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_88 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_89 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_90 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_92 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_93 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_94 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_95 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_97 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_98 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_99 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_100 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_101 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_102 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_103 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_104 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_105 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_106 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_107 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_108 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_109 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_13 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_36 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_34 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_117 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_118 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_119 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_121 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_123 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_126 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_127 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_122 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_124 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_120 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_125 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_128 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_129 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_130 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_131 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_132 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_134 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_135 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_136 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_137 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_138 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_139 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_140 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_141 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_142 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_143 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_144 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_145 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_146 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_147 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_148 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_149 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_150 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_151 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_152 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_154 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_155 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_156 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_157 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_158 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_159 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_160 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_161 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_162 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_163 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_164 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_165 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_166 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_167 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_168 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_169 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_170 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_171 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_172 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_173 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_174 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_175 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_176 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_177 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_178 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_179 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_180 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_181 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_183 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_182 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_184 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_186 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_187 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_188 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_189 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_190 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_191 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_192 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_193 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_194 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_195 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_196 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_197 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_198 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_199 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_200 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_201 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_202 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_203 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_204 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_205 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_206 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_207 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_208 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_209 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_210 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_211 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_212 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_213 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_214 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_215 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_216 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_217 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_218 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_219 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_220 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_221 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_222 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_223 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_224 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_225 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_226 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_227 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_228 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_229 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_230 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_231 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_232 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_233 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_247 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_248 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_249 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_250 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_251 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_252 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_253 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_265 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_275 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_274 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_273 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_272 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_271 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_11 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_12 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_13 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_14 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_15 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_16 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_17 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_18 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_19 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_20 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_21 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_22 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_286 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_287 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_288 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_289 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_290 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_23 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_24 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_25 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_26 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_27 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_28 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_29 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_30 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_31 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_32 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_33 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_34 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_35 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_36 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_37 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_38 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_39 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_40 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_41 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_42 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_43 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_44 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_45 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_46 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_47 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_48 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_49 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_50 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_51 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_52 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_53 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_54 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_55 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_56 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_57 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_58 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_59 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_60 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_61 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_62 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_64 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_67 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_68 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_69 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_71 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_72 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_73 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_74 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_75 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_76 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_77 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_78 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_79 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_80 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_81 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_82 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_83 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_84 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_85 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_87 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_88 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_89 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_90 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_92 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_93 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_95 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_96 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_97 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_98 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_99 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_101 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_102 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_104 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_105 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_107 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_108 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_109 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_110 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_112 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_113 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_114 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_115 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_117 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_118 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_119 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_120 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_121 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_122 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_123 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_125 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_126 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_127 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_129 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_130 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_131 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_132 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_134 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_135 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_136 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_138 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_139 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_140 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_142 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_143 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_144 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_146 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_148 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_149 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_150 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_151 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_153 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_154 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_155 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_156 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_157 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_159 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_161 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_162 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_163 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_164 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_165 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_167 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_169 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_170 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_171 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_172 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_173 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_174 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_175 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_176 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_177 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_179 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_180 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_182 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_291 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_300 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_10 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_183 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_184 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_185 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_186 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_187 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_188 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_189 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_190 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_191 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_192 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_193 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_270 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_194 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_195 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_196 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_197 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_198 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_199 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_200 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_201 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_202 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_203 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_204 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_205 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_206 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_207 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_208 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_209 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_210 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_211 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_212 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_213 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_215 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_214 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_216 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_217 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_218 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_219 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_220 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_221 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_222 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_223 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_224 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_225 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_226 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_227 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_228 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_229 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_230 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_231 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_232 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_233 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_234 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_235 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_236 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_237 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_238 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_239 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_240 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_241 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_242 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_243 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_244 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_245 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_246 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_247 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_248 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_185 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_249 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_269 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_250 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_251 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_252 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_253 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_254 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_255 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_256 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_257 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_258 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_259 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_260 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_261 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_262 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_263 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_264 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_265 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_266 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_267 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_268 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_269 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_270 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_271 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_272 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_273 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_274 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_275 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_276 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_277 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_278 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_279 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_280 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_281 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_282 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_283 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_284 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_285 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_286 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_287 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_288 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_289 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_290 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_291 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_292 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_268 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_293 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_294 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_267 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_302 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_303 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_295 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_296 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_306 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_307 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_308 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_309 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_310 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_311 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_312 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_313 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_314 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_266 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_315 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_316 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_317 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_318 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_319 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_320 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_321 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_322 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_323 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_324 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_325 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_326 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_327 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_328 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_329 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_330 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_331 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_332 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_336 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_337 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_338 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_341 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_342 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_343 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_344 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_347 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_351 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_352 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_353 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_356 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_360 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_361 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_362 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_365 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_369 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_370 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_371 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_374 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_378 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_379 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_382 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_386 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_285 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_422 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_423 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_424 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_284 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_425 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_446 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_447 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_448 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_449 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_450 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_451 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_452 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_453 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_283 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_23 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_282 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_281 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_280 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_21 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_81 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_78 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_279 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_278 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_277 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_276 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_39 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_40 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_32 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_28 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_29 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_33 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_48 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_51 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_56 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_57 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_14 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_363 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_364 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_366 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_389 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_466 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_392 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_390 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_393 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_467 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_394 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_468 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_472 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_473 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_297 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_298 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xana_filler_234 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_235 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_236 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_237 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_238 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_239 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_240 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_241 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_242 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_243 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_244 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_245 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_246 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_254 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_255 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xana_filler_256 TI1L1ASP10C1K2 $PINS AVSS=GNDD_IN AVDD=VDDH_IN 
Xd_fill_cap_178 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_181 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_299 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_300 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_301 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_302 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_303 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_304 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_305 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_333 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_334 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_335 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_339 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
Xd_fill_cap_340 TI1L1SP10C1K $PINS VSS=GNDD_IN VDD3=VDDH_IN 
