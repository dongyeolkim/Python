
*.BIPOLAR
*.RESVAL
*.CAPVAL

*.CONNECT VCC VCCNW
* TECHNOLOGY: FOF0L_PRS25
* CELL NAME : XOSCHINTLA
* FILE: NETLIST.LUMPED
* CREATED: TUE APR 15 15:01:33 2014
* PROGRAM "CALIBRE *XRC"
* VERSION "V2011.1_49.39"
* 
*.GLOBAL VCC2I  VCC2O  VCC2IO  VCC3I  VCC3O  VCC3IO  VCC18I  VCC18O  VCC18IO  VCC1I 
*+ VCC1O  VCC12I  VCC12O  VCC12IO  VCCK  VCCNW  VCC12A  VCC10A  VCC2A  VCC3A  VCC15IO 
*+ GND  GNDK  GNDI  GNDB  GNDO  GNDIO  GNDA  VCC 
.SUBCKT XOSCHINTLA O I IO E EB S0 S1 FEB
*XRI2335 N_1 VCC3IO VCC3IO RNPD_LP RN=49251.4 W=5E-07 L=0.0001435 
MI589 GNDIO N_1 GNDIO GNDIO N_25OD33_LP L=2.69E-05 W=2.9685E-05
MI2326 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_2 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2328 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2326-_2 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_3 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_4 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2326-_3 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_5 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_6 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2328-_2 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2328-_3 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2326-_4 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_7 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_8 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2326-_5 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_9 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_10 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2328-_4 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2328-_5 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2326-_6 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_11 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_12 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2326-_7 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_13 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_14 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2328-_6 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2326-_8 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_15 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_16 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2328-_7 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2326-_9 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_17 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_18 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2328-_8 N_2 N_1 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI2326-_10 VCC3IO N_2 GNDIO GNDIO N_25OD33_LP L=5E-07 W=4.1E-05
MI2327-_19 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI2327-_20 VCC3IO N_2 GNDK GNDK N_25OD33_LP L=5E-07 W=2.748E-05
MI590 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_2 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_3 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_4 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_5 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_6 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_7 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_8 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_9 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_10 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_11 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI590-_12 VCC3IO N_1 N_2 VCC3IO P_25OD33_LP L=4.2E-07 W=1.2E-05
MI_265 VCC3IO N_18 N_23 VCC3IO P_25OD33_LP L=4.2E-07 W=6E-06
MI_265-_2 VCC3IO N_18 N_23 VCC3IO P_25OD33_LP L=4.2E-07 W=6E-06
MI4626 VCC3IO VCC3IO N_69 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI_329 VCC3IO N_25 N_69 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
*XDI4688-_2 IO VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4688 IO VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4630-_2 I VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4630-_3 I VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4630-_4 I VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4630-_5 I VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4630 I VCC3IO DIOP_25_LP  AREA=1.4567E-10 PJ=0.00014042
*XDI4687-_2 GNDIO IO DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XDI4687 GNDIO IO DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XDI4629-_2 GNDIO I DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XDI4629-_3 GNDIO I DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XDI4629-_4 GNDIO I DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XDI4629-_5 GNDIO I DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XDI4629 GNDIO I DION_25_LP  AREA=9.36678E-11 PJ=9.182E-05
*XRI4681 IO N_68 VCC3IO RNPPO_LP RN=73.3054 W=7.45E-06 L=7E-07 
*XRI4682 IO N_26 VCC3IO RNPPO_LP RN=73.3054 W=7.45E-06 L=7E-07 
*XRI4679 IO N_22 VCC3IO RNPPO_LP RN=73.3054 W=7.45E-06 L=7E-07 
*XRI4678 IO N_23 VCC3IO RNPPO_LP RN=347.147 W=3.3E-06 L=1.52E-06 
*XRI4680 IO N_69 VCC3IO RNPPO_LP RN=73.3054 W=7.45E-06 L=7E-07 
MI_262 N_23 N_21 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI_262-_2 N_23 N_21 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI_324 N_69 N_24 GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI4623 N_69 GNDIO GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI4624 N_68 GNDIO GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI4622 N_68 N_24 GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI_55 N_26 N_20 GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI2105 N_26 GNDIO GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI2587 N_22 GNDIO GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI_211 N_22 N_17 GNDIO GNDIO N_25OD33_LP L=5E-07 W=2.93E-05
MI4626-_2 VCC3IO VCC3IO N_69 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI4627 VCC3IO VCC3IO N_68 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI4627-_2 VCC3IO VCC3IO N_68 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI2588 VCC3IO EPU N_26 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI2588-_2 VCC3IO EPU N_26 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI2589 VCC3IO VCC3IO N_22 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI2589-_2 VCC3IO VCC3IO N_22 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI_329-_2 VCC3IO N_25 N_69 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI4625 VCC3IO N_25 N_68 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI4625-_2 VCC3IO N_25 N_68 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI_56 VCC3IO N_19 N_26 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI_56-_2 VCC3IO N_19 N_26 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI_216 VCC3IO N_16 N_22 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
MI_216-_2 VCC3IO N_16 N_22 VCC3IO P_25OD33_LP L=4.2E-07 W=3.25E-05
*XRI710 N_66 I VCC3IO RNPPO_LP RN=345.923 W=2.6E-06 L=1.18E-06 
MI2349 EB3 ENG N_5 GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2254 ENG ENGB GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2348 N_5 S0S GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2347 GNDIO S1S N_5 GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2291 GPR GNR GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2202 N_57 TIEVC N_23 GNDK N_25OD33_LP L=5E-07 W=5E-06
MI2138 N_21 EB1 GNDIO GNDK N_25OD33_LP L=5E-07 W=2E-06
MI2202-_2 N_57 TIEVC N_23 GNDK N_25OD33_LP L=5E-07 W=5E-06
MI2139 N_17 EB3 GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2220 N_40 GNR N_57 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2221 N_41 GNR N_40 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2222 N_42 GNR N_41 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2223 N_43 GNR N_42 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2216 N_44 GNR N_43 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2217 N_45 GNR N_44 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2218 N_46 GNR N_45 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2219 N_47 GNR N_46 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2224 N_48 GNR N_47 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2225 N_49 GNR N_48 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2226 N_50 GNR N_49 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2227 N_51 GNR N_50 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2228 N_52 GNR N_51 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI_403 N_67 GNR N_52 GNDK N_25OD33_LP L=1.3E-05 W=7E-07
MI2255 EPU N_9 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2262 EEB N_11 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2261 _EEB EEB VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2286 GPR GNR VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2286-_2 GPR GNR VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2305 N_30 N_33 N_29 VCC3IO P_25OD33_LP L=4.2E-07 W=8E-07
MI2298 N_23 TIEGND N_57 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2298-_2 N_23 TIEGND N_57 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2207 N_57 GPR N_40 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2208 N_40 GPR N_41 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2209 N_41 GPR N_42 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2210 N_42 GPR N_43 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2203 N_43 GPR N_44 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2204 N_44 GPR N_45 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2205 N_45 GPR N_46 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2206 N_46 GPR N_47 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2211 N_47 GPR N_48 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2212 N_48 GPR N_49 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2213 N_49 GPR N_50 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2214 N_50 GPR N_51 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI2215 N_51 GPR N_52 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI_435 N_52 GPR N_67 VCC3IO P_25OD33_LP L=6E-06 W=7E-07
MI4247 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI4247-_2 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI4247-_3 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI4247-_4 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI2146 N_67 EB6 N_20 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2146-_2 N_67 EB6 N_20 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2144 N_67 EB6 N_19 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2144-_2 N_67 EB6 N_19 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2147 N_67 EB8 N_24 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2147-_2 N_67 EB8 N_24 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2148 N_67 EB8 N_25 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2148-_2 N_67 EB8 N_25 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2306 N_33 N_27 N_29 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2307 N_29 N_27 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2302 N_20 EB5 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2302-_2 N_20 EB5 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2303 N_19 EB5 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2303-_2 N_19 EB5 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2300 N_24 EB7 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2300-_2 N_24 EB7 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2301 N_25 EB7 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2301-_2 N_25 EB7 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2304 N_31 TIEGND VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=3E-06
MI2330 VCC3IO N_62 N_62 VCC3IO P_25OD33_LP L=4.2E-07 W=3E-06
MI_127 N_19 EB6 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=3E-06
MI_127-_2 N_19 EB6 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=3E-06
MI_328 N_25 EB8 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=3E-06
MI_328-_2 N_25 EB8 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=3E-06
MI_193 N_30 TIEVC GNDIO GNDK N_25OD33_LP L=5E-07 W=3E-06
MI2145 N_20 EB5 GNDIO GNDK N_25OD33_LP L=5E-07 W=3E-06
MI_325 N_24 EB7 GNDIO GNDK N_25OD33_LP L=5E-07 W=3E-06
MI2141 N_67 EB2 N_21 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2140 N_67 EB2 N_18 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2143 N_67 EB4 N_17 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2142 N_67 EB4 N_16 GNDK N_25OD33_LP L=5E-07 W=2.5E-06
MI2317 N_21 EB1 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2318 N_18 EB1 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2315 N_17 EB3 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2314 N_16 EB3 N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2321 N_32 N_33 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI4677 N_70 N_32 VCCK VCCK P_25OD33_LP L=4.2E-07 W=2E-06
MI4677-_2 N_70 N_32 VCCK VCCK P_25OD33_LP L=4.2E-07 W=2E-06
MI_264 N_18 EB2 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI_215 N_16 EB4 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI2137 N_57 EEB N_27 GNDK N_25OD33_LP L=5E-07 W=1.25E-06
MI2137-_2 N_57 EEB N_27 GNDK N_25OD33_LP L=5E-07 W=1.25E-06
MI2299 N_27 _EEB N_57 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2299-_2 N_27 _EEB N_57 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-06
MI2329 TIEGND N_62 GNDIO GNDK N_25OD33_LP L=5E-07 W=4E-06
MI2331 N_61 N_61 GNDIO GNDK N_25OD33_LP L=5E-07 W=4E-06
MI2331-_2 N_61 N_61 GNDIO GNDK N_25OD33_LP L=5E-07 W=4E-06
MI2332 VCC3IO N_61 TIEVC VCC3IO P_25OD33_LP L=4.2E-07 W=4E-06
MI2332-_2 VCC3IO N_61 TIEVC VCC3IO P_25OD33_LP L=4.2E-07 W=4E-06
MI4248 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_2 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_3 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_4 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_5 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_6 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_7 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI4248-_8 O N_70 GNDK GNDK N_12_LPRVT L=6E-08 W=5E-07
MI_194 N_31 N_33 N_28 GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2136 N_27 _EEB GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI4676 N_70 N_32 GNDK GNDK N_25OD33_LP L=5E-07 W=1E-06
MI4676-_2 N_70 N_32 GNDK GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2323 N_32 N_33 GNDIO GNDK N_25OD33_LP L=5E-07 W=2E-06
MI2323-_2 N_32 N_33 GNDIO GNDK N_25OD33_LP L=5E-07 W=2E-06
MI4247-_5 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI4247-_6 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI4247-_7 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI4247-_8 VCCK N_70 O VCCK P_12_LPRVT L=6E-08 W=1E-06
MI_195 N_33 N_27 N_28 GNDK N_25OD33_LP L=5E-07 W=2.7E-06
MI2118 N_28 N_27 GNDIO GNDK N_25OD33_LP L=5E-07 W=2.7E-06
*XDI4637 GNDK E DION_12_LPRVT  AREA=1.421E-13 PJ=1.56E-06
*XDI4686 GNDK EB DION_12_LPRVT  AREA=1.421E-13 PJ=1.56E-06
*XDI4683 GNDK FEB DION_12_LPRVT  AREA=1.421E-13 PJ=1.56E-06
*XDI4684 GNDK S0 DION_12_LPRVT  AREA=1.421E-13 PJ=1.56E-06
*XDI4685 GNDK S1 DION_12_LPRVT  AREA=1.421E-13 PJ=1.56E-06
MI2253 N_15 _EB2V GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2252 ENGB E2V N_15 GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2259 N_9 E2V GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2258 EPU N_9 GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2260 N_9 EB2V GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2266 EEB N_11 GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2267 N_11 E2V GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2265 _EEB EEB GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2268 N_11 _EB2V GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2292 GNR FEB2V GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI2293 GNR ENGB GNDIO GNDK N_25OD33_LP L=5E-07 W=7E-07
MI4639 VCCK E N_36 VCCK P_12_LPRVT L=6E-08 W=5E-07
MI4638 N_36 E GNDK GNDK N_12_LPRVT L=6E-08 W=3E-07
MI4632 E2V N_36 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4631 _E2V E GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4636 VCC3IO _E2V N_35 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4633 N_35 N_36 E2V VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4634 VCC3IO E2V N_34 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4635 N_34 E _E2V VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4648 VCCK EB N_39 VCCK P_12_LPRVT L=6E-08 W=5E-07
MI4647 N_39 EB GNDK GNDK N_12_LPRVT L=6E-08 W=3E-07
MI4641 EB2V N_39 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4640 _EB2V EB GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4645 VCC3IO _EB2V N_38 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4642 N_38 N_39 EB2V VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4643 VCC3IO EB2V N_37 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4644 N_37 EB _EB2V VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4657 VCCK FEB N_56 VCCK P_12_LPRVT L=6E-08 W=5E-07
MI4656 N_56 FEB GNDK GNDK N_12_LPRVT L=6E-08 W=3E-07
MI4650 FEB2V N_56 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4649 N_53 FEB GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4654 VCC3IO N_53 N_55 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4651 N_55 N_56 FEB2V VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4652 VCC3IO FEB2V N_54 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4653 N_54 FEB N_53 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4675 VCCK S0 N_60 VCCK P_12_LPRVT L=6E-08 W=5E-07
MI4673 N_60 S0 GNDK GNDK N_12_LPRVT L=6E-08 W=3E-07
MI4661 S0S N_60 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4660 S0B S0 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4669 VCC3IO S0B N_59 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4666 N_59 N_60 S0S VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4667 VCC3IO S0S N_58 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4668 N_58 S0 S0B VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4674 VCCK S1 N_65 VCCK P_12_LPRVT L=6E-08 W=5E-07
MI4672 N_65 S1 GNDK GNDK N_12_LPRVT L=6E-08 W=3E-07
MI4659 S1S N_65 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4658 S1B S1 GNDK GNDK N_25OD33_LP L=5E-07 W=8.8E-06
MI4665 VCC3IO S1B N_64 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4662 N_64 N_65 S1S VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4664 VCC3IO S1S N_63 VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI4663 N_63 S1 S1B VCC3IO P_25OD33_LP L=4.2E-07 W=5E-07
MI2256 N_9 EB2V N_8 VCC3IO P_25OD33_LP L=4.2E-07 W=1.4E-06
MI2263 N_11 _EB2V N_10 VCC3IO P_25OD33_LP L=4.2E-07 W=1.4E-06
MI2287 GNR ENGB N_7 VCC3IO P_25OD33_LP L=4.2E-07 W=1.4E-06
MI2257 N_8 E2V VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1.4E-06
MI2264 N_10 E2V VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1.4E-06
MI2288 N_7 FEB2V VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1.4E-06
MI2346 EB4 EB3 GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2341 EB1 ENG GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2340 EB2 EB1 GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2192 N_12 S0S GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2174 EB6 EB5 GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2193 EB5 ENG N_12 GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2190 EB7 ENG N_13 GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2173 EB8 EB7 GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2189 N_13 S0S N_14 GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2188 N_14 S1S GNDIO GNDK N_25OD33_LP L=5E-07 W=1E-06
MI2250 ENGB _EB2V VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2251 ENG ENGB VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2343 EB3 ENG VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2249 ENGB E2V VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2339 EB1 ENG VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2345 VCC3IO S0S N_6 VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2344 N_6 S1S EB3 VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2181 EB5 S0S VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2182 EB5 ENG VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2179 EB7 ENG VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2178 EB7 S0S VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2177 EB7 S1S VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=1E-06
MI2342 EB4 EB3 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI2338 EB2 EB1 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI2170 EB6 EB5 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI2169 EB8 EB7 VCC3IO VCC3IO P_25OD33_LP L=4.2E-07 W=2E-06
MI2334 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_2 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_3 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_4 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_5 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_6 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_7 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_8 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_9 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_10 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_11 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_12 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_13 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_14 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_15 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=5E-06
MI2334-_16 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_17 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_18 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_19 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_20 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_21 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2334-_22 VCC3IO GNDIO VCC3IO VCC3IO P_25OD33_LP L=5E-06 W=1E-05
MI2200 N_67 TIEVC N_66 GNDK N_25OD33_LP L=5E-07 W=7.5E-06
MI2200-_2 N_67 TIEVC N_66 GNDK N_25OD33_LP L=5E-07 W=7.5E-06
MI2316 N_66 TIEGND N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=7.5E-06
MI2316-_2 N_66 TIEGND N_67 VCC3IO P_25OD33_LP L=4.2E-07 W=7.5E-06
*XRI2336 N_4 VCCK VCCK RNPD_LP RN=49251.4 W=5E-07 L=0.0001435 
MI2333 GNDIO N_4 GNDIO GNDIO N_25OD33_LP L=2.69E-05 W=2.9685E-05
MI587 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_2 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_3 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_4 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_5 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_6 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_7 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI587-_8 N_3 N_4 GNDIO GNDIO N_25OD33_LP L=5E-07 W=3E-06
MI405 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_2 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_3 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_4 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_5 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_6 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_7 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_8 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_9 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_10 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_11 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI405-_12 VCCK N_4 N_3 VCCK P_25OD33_LP L=4.2E-07 W=1.2E-05
MI588 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI588-_2 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_3 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_4 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI588-_5 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_6 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_7 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI588-_8 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_9 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_10 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI588-_11 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_12 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_13 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI588-_14 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI588-_15 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI399-_2 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_3 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_4 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI399-_5 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_6 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_7 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI399-_8 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_9 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_10 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI399-_11 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_12 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_13 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=4.1E-05
MI399-_14 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
MI399-_15 VCCK N_3 GNDIO GNDIO N_12_LPRVT L=9E-08 W=2.748E-05
*.ENDS
*
*
.SUBCKT P_12_LPLVT D G S B W=W L=L
M0 D G S B P_12_LPLVT W=W L=L
.ENDS

.SUBCKT P_12_LPRVT D G S B W=W L=L
M1 D G S B P_12_LPRVT W=W L=L
.ENDS

.SUBCKT P_12_LPHVT D G S B W=W L=L
M1 D G S B P_12_LPHVT W=W L=L
.ENDS

.SUBCKT P_25_LP D G S B W=W L=L
M1 D G S B P_25_LP W=W L=L
.ENDS

.SUBCKT P_25OD33_LP D G S B W=W L=L
M1 D G S B P_25OD33_LP W=W L=L
.ENDS

.SUBCKT P_25UD18_LP D G S B W=W L=L
M1 D G S B P_25UD18_LP W=W L=L
.ENDS

.SUBCKT P_L42P5_LPHVT D G S B W=W L=L
M1 D G S B P_L42P5_LPHVT W=W L=L
.ENDS

.SUBCKT P_L52P5_ULPHVT D G S B W=W L=L
M1 D G S B P_L52P5_ULPHVT W=W L=L
.ENDS

.SUBCKT P_L78P9_LPHVT D G S B W=W L=L
M1 D G S B P_L78P9_LPHVT W=W L=L
.ENDS

.SUBCKT N_12_LPLVT D G S B W=W L=L
M0 D G S B N_12_LPLVT W=W L=L
.ENDS

.SUBCKT N_BPW_12_LPLVT D G S B W=W L=L
M0 D G S B N_BPW_12_LPLVT W=W L=L
.ENDS

.SUBCKT N_BPW_12_LPRVT D G S B W=W L=L
M1 D G S B N_BPW_12_LPRVT W=W L=L
.ENDS

.SUBCKT N_12_LPRVT D G S B W=W L=L
M1 D G S B N_12_LPRVT W=W L=L
.ENDS

.SUBCKT N_BPW_12_LPHVT W=W L=L
M1 D G S B N_BPW_12_LPHVT W=W L=L
.ENDS

.SUBCKT N_12_LPHVT D G S B W=W L=L
M1 D G S B N_12_LPHVT W=W L=L
.ENDS

.SUBCKT N_12_LPNVT D G S B W=W L=L
M1 D G S B N_12_LPNVT W=W L=L
.ENDS

.SUBCKT N_25_LP D G S B W=W L=L
M1 D G S B N_25_LP W=W L=L
.ENDS

.SUBCKT N_BPW_25_LP D G S B W=W L=L
M1 D G S B N_BPW_25_LP W=W L=L
.ENDS

.SUBCKT N_25OD33_LP D G S B W=W L=L
M1 D G S B N_25OD33_LP W=W L=L
.ENDS

.SUBCKT N_BPW_25OD33_LP D G S B W=W L=L
M1 D G S B N_BPW_25OD33_LP W=W L=L
.ENDS

.SUBCKT RNNPO_LP POS NEG SUB
R0 POS NEG RNNPO_LP R=RN $SUB=SUB
.ENDS

.SUBCKT RNPPO_LP POS NEG WEL
R1 POS NEG RNPPO_LP R=RN $SUB=WEL
.ENDS

.SUBCKT RNND_LP POS NEG SUB
R0 POS NEG RNND_LP R=RN $SUB=SUB
.ENDS

.SUBCKT RNPD_LP POS NEG WEL
R1 POS NEG RNPD_LP R=RN $SUB=WEL
.ENDS

.SUBCKT RSNWELP_LP POS NEG SUB
R0 POS NEG RSNWELP_LP R=RN $SUB=SUB
.ENDS

.SUBCKT RSND_LP POS NEG SUB
R0 POS NEG RSND_LP R=RN $SUB=SUB
.ENDS

.SUBCKT RSPD_LP POS NEG WEL
R0 POS NEG RSPD_LP R=RN $SUB=WEL
.ENDS

.SUBCKT RSNPO_LP POS NEG SUB
R0 POS NEG RSNPO_LP R=RN $SUB=SUB
.ENDS

.SUBCKT RSPPO_LP POS NEG WEL
R0 POS NEG RSPPO_LP R=RN $SUB=WEL
.ENDS

.SUBCKT RSNWELL_LP POS NEG SUB
R0 POS NEG RSNWELL_LP R=RN $SUB=SUB
.ENDS

.SUBCKT DIOP_12_LPRVT POS NEG AREA=AREA PJ=PJ
D0 POS NEG DIOP_12_LPRVT AREA=AREA PJ=PJ
.ENDS

.SUBCKT DIOP_12_LPHVT POS NEG AREA=AREA PJ=PJ
D0 POS NEG DIOP_12_LPHVT AREA=AREA PJ=PJ
.ENDS

.SUBCKT DIOP_12_LPLVT POS NEG AREA=AREA PJ=PJ
D0 POS NEG DIOP_12_LPLVT AREA=AREA PJ=PJ
.ENDS

.SUBCKT DION_12_LPRVT POS NEG AREA=AREA PJ=PJ
D0 POS NEG DION_12_LPRVT AREA=AREA PJ=PJ
.ENDS

.SUBCKT DION_12_LPHVT POS NEG AREA=AREA PJ=PJ
D0 POS NEG DION_12_LPHVT AREA=AREA PJ=PJ
.ENDS

.SUBCKT DION_12_LPLVT POS NEG AREA=AREA PJ=PJ
D0 POS NEG DION_12_LPLVT AREA=AREA PJ=PJ
.ENDS

.SUBCKT DIOP_25_LP POS NEG AREA=AREA PJ=PJ
D0 POS NEG DIOP_25_LP AREA=AREA PJ=PJ
.ENDS

.SUBCKT DION_25_LP POS NEG AREA=AREA PJ=PJ
D0 POS NEG DION_25_LP AREA=AREA PJ=PJ
.ENDS

.SUBCKT DIONW_25_LP POS NEG AREA=AREA PJ=PJ
D0 POS NEG DIONW_25_LP AREA=AREA PJ=PJ
.ENDS

.SUBCKT NCAP_12_LP POS NEG
C0 POS NEG NCAP_12_LP NF=NF WF=WF LF=LF
.ENDS

.SUBCKT NCAP_25_LP POS NEG
C0 POS NEG NCAP_25_LP NF=NF WF=WF LF=LF
.ENDS

.SUBCKT NCAP_33_LP POS NEG
C0 POS NEG NCAP_33_LP NF=NF WF=WF LF=LF
.ENDS

.SUBCKT P_12_ULPUHVT D G S B W=W L=L
M1 D G S B P_12_ULPUHVT W=W L=L
.ENDS

.SUBCKT N_12_ULPUHVT D G S B W=W L=L
M1 D G S B N_12_ULPUHVT W=W L=L
.ENDS

.end
